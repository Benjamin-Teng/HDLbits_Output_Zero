module moduleName (
    output zero
);
    
endmodule